magic
tech sky130A
timestamp 1763960441
<< nwell >>
rect -145 90 90 240
<< nmos >>
rect -5 -50 10 50
<< pmos >>
rect -5 115 10 215
<< ndiff >>
rect -65 35 -5 50
rect -65 -35 -50 35
rect -20 -35 -5 35
rect -65 -50 -5 -35
rect 10 35 70 50
rect 10 -35 25 35
rect 55 -35 70 35
rect 10 -50 70 -35
<< pdiff >>
rect -65 200 -5 215
rect -65 130 -50 200
rect -20 130 -5 200
rect -65 115 -5 130
rect 10 200 70 215
rect 10 130 25 200
rect 55 130 70 200
rect 10 115 70 130
<< ndiffc >>
rect -50 -35 -20 35
rect 25 -35 55 35
<< pdiffc >>
rect -50 130 -20 200
rect 25 130 55 200
<< psubdiff >>
rect -125 35 -65 50
rect -125 -35 -110 35
rect -80 -35 -65 35
rect -125 -50 -65 -35
<< nsubdiff >>
rect -125 200 -65 215
rect -125 130 -110 200
rect -80 130 -65 200
rect -125 115 -65 130
<< psubdiffcont >>
rect -110 -35 -80 35
<< nsubdiffcont >>
rect -110 130 -80 200
<< poly >>
rect -5 215 10 230
rect -5 50 10 115
rect -5 -70 10 -50
rect -45 -80 10 -70
rect -45 -100 -35 -80
rect -15 -85 10 -80
rect -15 -100 -5 -85
rect -45 -110 -5 -100
<< polycont >>
rect -35 -100 -15 -80
<< locali >>
rect -120 200 -10 210
rect -120 130 -110 200
rect -80 130 -50 200
rect -20 130 -10 200
rect -120 120 -10 130
rect 15 200 65 210
rect 15 130 25 200
rect 55 130 65 200
rect 15 120 65 130
rect 25 45 55 120
rect -120 35 -10 45
rect -120 -35 -110 35
rect -80 -35 -50 35
rect -20 -35 -10 35
rect -120 -45 -10 -35
rect 15 35 65 45
rect 15 -35 25 35
rect 55 -35 65 35
rect 15 -45 65 -35
rect 25 -65 55 -45
rect -145 -80 -5 -75
rect -145 -100 -35 -80
rect -15 -100 -5 -80
rect 25 -90 70 -65
rect -145 -105 -5 -100
<< viali >>
rect -110 130 -80 200
rect -50 130 -20 200
rect -110 -35 -80 35
rect -50 -35 -20 35
<< metal1 >>
rect -145 200 -10 210
rect -145 130 -110 200
rect -80 130 -50 200
rect -20 130 -10 200
rect -145 120 -10 130
rect -145 35 -10 45
rect -145 -35 -110 35
rect -80 -35 -50 35
rect -20 -35 -10 35
rect -145 -45 -10 -35
<< labels >>
rlabel metal1 -145 165 -145 165 7 VDD
port 1 w
rlabel metal1 -145 0 -145 0 7 VSS
port 2 w
rlabel locali -145 -90 -145 -90 7 A
port 3 w
rlabel locali 70 -75 70 -75 3 Y
port 4 e
<< end >>
